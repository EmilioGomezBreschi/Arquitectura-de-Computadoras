
`timescale 1ns/1ns
 //definicion del modulo
module expresso(
    input [3:0]a,
    input [3:0]b,
    output [3:0]c
);
 //definicion de cables o registros 

 //cuerpo del modulo assigns(si) instancias(n/a) always(n/a)
    assign c = a + b; //se suma todo el rango de a con el de b, no se especifican bits


 endmodule