//inicio de modulo con inputs y outputs
module S32C(
	input [31:0]A,
	input [31:0]B,
	output [31:0]C
);

// asignaciones

assign C=A+B;

endmodule
